library verilog;
use verilog.vl_types.all;
entity CounterDown4_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end CounterDown4_vlg_sample_tst;
