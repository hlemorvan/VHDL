library verilog;
use verilog.vl_types.all;
entity RegisterN_vlg_vec_tst is
end RegisterN_vlg_vec_tst;
