library verilog;
use verilog.vl_types.all;
entity FlipFlopD_vlg_vec_tst is
end FlipFlopD_vlg_vec_tst;
