library verilog;
use verilog.vl_types.all;
entity CounterDown4_vlg_vec_tst is
end CounterDown4_vlg_vec_tst;
